`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:19:06 10/24/2016 
// Design Name: 
// Module Name:    ALU_Execute 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ALU_Execute(
   input [10:0] ctrl,
   input clk,
   input [5:0] reg1,
   input [5:0] reg2,
   input [63:0] se,
   input [3:0] aluCtrl
   );
	
	

endmodule
